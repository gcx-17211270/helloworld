//�߳��� 2020.04.20
//�������ķ��漤����
//testbench		tb

module inv_tb();

endmodule