//�߳���	2020.04.20
//����һ��������

module();



endmodule